module a0;
	int x, y, z;
	assign z = x - y - 1;
endmodule
