(* dont_touch = "true" *)
