entity foo is
end;

architecture bar of foo is
begin
end;

-- entity @foo_bar () () {
-- }
