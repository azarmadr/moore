// RUN: moore %s
module foo;
  int a;
  int b = a;
endmodule
