entity foo is end;
architecture bar of foo is
	constant TOLER: DISTANCE := 1.5 nm;
	constant PI: REAL := 3.141592;
	constant CYCLE_TIME: TIME := 100 ns;
	constant Propagation_Delay: DELAY_LENGTH;
begin end;
